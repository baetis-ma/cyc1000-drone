
module pll (
	clk_clk,
	reset_reset_n,
	pll_clk);	

	input		clk_clk;
	input		reset_reset_n;
	output		pll_clk;
endmodule
